module quicksort

pub fn sort[T](mut array []T) {
	
}
